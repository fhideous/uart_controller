`timescale 1ns / 1ps

module uart_allocation_tb;
    
    reg      clk;
    reg      reset;

    reg      rx_i;
    wire     tx_o;
    
    localparam CLK_SEMIPERIOD = 5;
    
uart_allocation uut
(

  .clk      (clk        ),
  .reset    (reset      ),

  .rx_i     (rx_i       ),
  .tx_o     (tx_o       )


);

  initial begin 
     clk = 'b0;
     forever begin
       #CLK_SEMIPERIOD clk = ~clk;
     end
  end

reg  [7:0]  data;

integer   CLKS_PER_BIT    = 100_000_000_0 / 9600;
 
 
 initial begin 


  reset = 'b0;
  rx_i = 1'b1;
  data = 8'b1;
 #5000;
  reset = 'b1;
 #5000;

  data = 8'b1000_0001;
      rx_i = 1'b1;
      #2000;

      //start bit
  rx_i = 1'b0;
  #CLKS_PER_BIT;
      //data
  rx_i = data[0];
  #CLKS_PER_BIT;
  rx_i = data[1];
  #CLKS_PER_BIT;
  rx_i = data[2];
  #CLKS_PER_BIT;
  rx_i = data[3];
  #CLKS_PER_BIT;
  rx_i = data[4];
  #CLKS_PER_BIT;
  rx_i = data[5];
  #CLKS_PER_BIT;
  rx_i = data[6];
  #CLKS_PER_BIT;
  rx_i = data[7];
  #CLKS_PER_BIT;
  // stop bit
  rx_i = 1'b1;
  #CLKS_PER_BIT;

  data = 8'b0010_0110;

      //start bit
  rx_i = 1'b0;
  #CLKS_PER_BIT;
      //data
  rx_i = data[0];
  #CLKS_PER_BIT;
  rx_i = data[1];
  #CLKS_PER_BIT;
  rx_i = data[2];
  #CLKS_PER_BIT;
  rx_i = data[3];
  #CLKS_PER_BIT;
  rx_i = data[4];
  #CLKS_PER_BIT;
  rx_i = data[5];
  #CLKS_PER_BIT;
  rx_i = data[6];
  #CLKS_PER_BIT;
  rx_i = data[7];
  #CLKS_PER_BIT;
  // stop bit
  rx_i = 1'b1;
  #CLKS_PER_BIT;

  #CLKS_PER_BIT;
  #CLKS_PER_BIT;
  #CLKS_PER_BIT;
  #CLKS_PER_BIT;
  #CLKS_PER_BIT;
  #CLKS_PER_BIT;
  #CLKS_PER_BIT;
  #CLKS_PER_BIT;
  #CLKS_PER_BIT;
  #CLKS_PER_BIT;
  #CLKS_PER_BIT;
  #CLKS_PER_BIT;
  #CLKS_PER_BIT;
  #CLKS_PER_BIT;
  #CLKS_PER_BIT;
  #CLKS_PER_BIT;
  #CLKS_PER_BIT;
  #CLKS_PER_BIT;
  #CLKS_PER_BIT;
  #CLKS_PER_BIT;

  data = 8'b1000_1000;

      //start bit
  rx_i = 1'b0;
  #CLKS_PER_BIT;
      //data
  rx_i = data[0];
  #CLKS_PER_BIT;
  rx_i = data[1];
  #CLKS_PER_BIT;
  rx_i = data[2];
  #CLKS_PER_BIT;
  rx_i = data[3];
  #CLKS_PER_BIT;
  rx_i = data[4];
  #CLKS_PER_BIT;
  rx_i = data[5];
  #CLKS_PER_BIT;
  rx_i = data[6];
  #CLKS_PER_BIT;
  rx_i = data[7];
  #CLKS_PER_BIT;
  // stop bit
  rx_i = 1'b1;
  #CLKS_PER_BIT;


 end




endmodule